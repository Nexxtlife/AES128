-- test_interface_sys.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity test_interface_sys is
	port (
		aes_interface_0_avalon_streaming_source_data  : out std_logic_vector(127 downto 0);        -- aes_interface_0_avalon_streaming_source.data
		aes_interface_0_avalon_streaming_source_ready : in  std_logic                      := '0'; --                                        .ready
		aes_interface_0_avalon_streaming_source_valid : out std_logic;                             --                                        .valid
		clk_clk                                       : in  std_logic                      := '0'; --                                     clk.clk
		reset_reset_n                                 : in  std_logic                      := '0'  --                                   reset.reset_n
	);
end entity test_interface_sys;

architecture rtl of test_interface_sys is
	component interface is
		port (
			interface_0_avalon_streaming_source_data  : out std_logic_vector(127 downto 0);                    -- data
			interface_0_avalon_streaming_source_ready : in  std_logic                      := 'X';             -- ready
			interface_0_avalon_streaming_source_valid : out std_logic;                                         -- valid
			clk_clk                                   : in  std_logic                      := 'X';             -- clk
			reset_reset_n                             : in  std_logic                      := 'X';             -- reset
			interface_0_avalon_master_1_address       : out std_logic_vector(16 downto 0);                     -- address
			interface_0_avalon_master_1_byteenable    : out std_logic_vector(15 downto 0);                     -- byteenable
			interface_0_avalon_master_1_read          : out std_logic;                                         -- read
			interface_0_avalon_master_1_readdata      : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			interface_0_avalon_master_1_waitrequest   : in  std_logic                      := 'X'              -- waitrequest
		);
	end component interface;

	component test_interface_sys_onchip_memory2_0 is
		port (
			clk         : in  std_logic                      := 'X';             -- clk
			address     : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			debugaccess : in  std_logic                      := 'X';             -- debugaccess
			clken       : in  std_logic                      := 'X';             -- clken
			chipselect  : in  std_logic                      := 'X';             -- chipselect
			write       : in  std_logic                      := 'X';             -- write
			readdata    : out std_logic_vector(127 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                      := 'X';             -- reset
			reset_req   : in  std_logic                      := 'X';             -- reset_req
			freeze      : in  std_logic                      := 'X'              -- freeze
		);
	end component test_interface_sys_onchip_memory2_0;

	component test_interface_sys_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                          : in  std_logic                      := 'X';             -- clk
			aes_interface_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			aes_interface_0_avalon_master_address                  : in  std_logic_vector(16 downto 0)  := (others => 'X'); -- address
			aes_interface_0_avalon_master_waitrequest              : out std_logic;                                         -- waitrequest
			aes_interface_0_avalon_master_byteenable               : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			aes_interface_0_avalon_master_read                     : in  std_logic                      := 'X';             -- read
			aes_interface_0_avalon_master_readdata                 : out std_logic_vector(127 downto 0);                    -- readdata
			onchip_memory2_0_s1_address                            : out std_logic_vector(2 downto 0);                      -- address
			onchip_memory2_0_s1_write                              : out std_logic;                                         -- write
			onchip_memory2_0_s1_readdata                           : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                          : out std_logic_vector(127 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                         : out std_logic_vector(15 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                         : out std_logic;                                         -- chipselect
			onchip_memory2_0_s1_clken                              : out std_logic;                                         -- clken
			onchip_memory2_0_s1_debugaccess                        : out std_logic                                          -- debugaccess
		);
	end component test_interface_sys_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal aes_interface_0_avalon_master_readdata            : std_logic_vector(127 downto 0); -- mm_interconnect_0:aes_interface_0_avalon_master_readdata -> aes_interface_0:interface_0_avalon_master_1_readdata
	signal aes_interface_0_avalon_master_waitrequest         : std_logic;                      -- mm_interconnect_0:aes_interface_0_avalon_master_waitrequest -> aes_interface_0:interface_0_avalon_master_1_waitrequest
	signal aes_interface_0_avalon_master_address             : std_logic_vector(16 downto 0);  -- aes_interface_0:interface_0_avalon_master_1_address -> mm_interconnect_0:aes_interface_0_avalon_master_address
	signal aes_interface_0_avalon_master_byteenable          : std_logic_vector(15 downto 0);  -- aes_interface_0:interface_0_avalon_master_1_byteenable -> mm_interconnect_0:aes_interface_0_avalon_master_byteenable
	signal aes_interface_0_avalon_master_read                : std_logic;                      -- aes_interface_0:interface_0_avalon_master_1_read -> mm_interconnect_0:aes_interface_0_avalon_master_read
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect  : std_logic;                      -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata    : std_logic_vector(127 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_debugaccess : std_logic;                      -- mm_interconnect_0:onchip_memory2_0_s1_debugaccess -> onchip_memory2_0:debugaccess
	signal mm_interconnect_0_onchip_memory2_0_s1_address     : std_logic_vector(2 downto 0);   -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable  : std_logic_vector(15 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write       : std_logic;                      -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata   : std_logic_vector(127 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken       : std_logic;                      -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal rst_controller_reset_out_reset                    : std_logic;                      -- rst_controller:reset_out -> [aes_interface_0:reset_reset_n, mm_interconnect_0:aes_interface_0_reset_sink_reset_bridge_in_reset_reset, onchip_memory2_0:reset]
	signal rst_controller_reset_out_reset_req                : std_logic;                      -- rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                           : std_logic;                      -- reset_reset_n:inv -> rst_controller:reset_in0

begin

	aes_interface_0 : component interface
		port map (
			interface_0_avalon_streaming_source_data  => aes_interface_0_avalon_streaming_source_data,  -- avalon_streaming_source.data
			interface_0_avalon_streaming_source_ready => aes_interface_0_avalon_streaming_source_ready, --                        .ready
			interface_0_avalon_streaming_source_valid => aes_interface_0_avalon_streaming_source_valid, --                        .valid
			clk_clk                                   => clk_clk,                                       --              clock_sink.clk
			reset_reset_n                             => rst_controller_reset_out_reset,                --              reset_sink.reset
			interface_0_avalon_master_1_address       => aes_interface_0_avalon_master_address,         --           avalon_master.address
			interface_0_avalon_master_1_byteenable    => aes_interface_0_avalon_master_byteenable,      --                        .byteenable
			interface_0_avalon_master_1_read          => aes_interface_0_avalon_master_read,            --                        .read
			interface_0_avalon_master_1_readdata      => aes_interface_0_avalon_master_readdata,        --                        .readdata
			interface_0_avalon_master_1_waitrequest   => aes_interface_0_avalon_master_waitrequest      --                        .waitrequest
		);

	onchip_memory2_0 : component test_interface_sys_onchip_memory2_0
		port map (
			clk         => clk_clk,                                           --   clk1.clk
			address     => mm_interconnect_0_onchip_memory2_0_s1_address,     --     s1.address
			debugaccess => mm_interconnect_0_onchip_memory2_0_s1_debugaccess, --       .debugaccess
			clken       => mm_interconnect_0_onchip_memory2_0_s1_clken,       --       .clken
			chipselect  => mm_interconnect_0_onchip_memory2_0_s1_chipselect,  --       .chipselect
			write       => mm_interconnect_0_onchip_memory2_0_s1_write,       --       .write
			readdata    => mm_interconnect_0_onchip_memory2_0_s1_readdata,    --       .readdata
			writedata   => mm_interconnect_0_onchip_memory2_0_s1_writedata,   --       .writedata
			byteenable  => mm_interconnect_0_onchip_memory2_0_s1_byteenable,  --       .byteenable
			reset       => rst_controller_reset_out_reset,                    -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,                --       .reset_req
			freeze      => '0'                                                -- (terminated)
		);

	mm_interconnect_0 : component test_interface_sys_mm_interconnect_0
		port map (
			clk_0_clk_clk                                          => clk_clk,                                           --                                        clk_0_clk.clk
			aes_interface_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                    -- aes_interface_0_reset_sink_reset_bridge_in_reset.reset
			aes_interface_0_avalon_master_address                  => aes_interface_0_avalon_master_address,             --                    aes_interface_0_avalon_master.address
			aes_interface_0_avalon_master_waitrequest              => aes_interface_0_avalon_master_waitrequest,         --                                                 .waitrequest
			aes_interface_0_avalon_master_byteenable               => aes_interface_0_avalon_master_byteenable,          --                                                 .byteenable
			aes_interface_0_avalon_master_read                     => aes_interface_0_avalon_master_read,                --                                                 .read
			aes_interface_0_avalon_master_readdata                 => aes_interface_0_avalon_master_readdata,            --                                                 .readdata
			onchip_memory2_0_s1_address                            => mm_interconnect_0_onchip_memory2_0_s1_address,     --                              onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                              => mm_interconnect_0_onchip_memory2_0_s1_write,       --                                                 .write
			onchip_memory2_0_s1_readdata                           => mm_interconnect_0_onchip_memory2_0_s1_readdata,    --                                                 .readdata
			onchip_memory2_0_s1_writedata                          => mm_interconnect_0_onchip_memory2_0_s1_writedata,   --                                                 .writedata
			onchip_memory2_0_s1_byteenable                         => mm_interconnect_0_onchip_memory2_0_s1_byteenable,  --                                                 .byteenable
			onchip_memory2_0_s1_chipselect                         => mm_interconnect_0_onchip_memory2_0_s1_chipselect,  --                                                 .chipselect
			onchip_memory2_0_s1_clken                              => mm_interconnect_0_onchip_memory2_0_s1_clken,       --                                                 .clken
			onchip_memory2_0_s1_debugaccess                        => mm_interconnect_0_onchip_memory2_0_s1_debugaccess  --                                                 .debugaccess
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of test_interface_sys
