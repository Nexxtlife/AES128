-- byteSub_display_sys.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity byteSub_display_sys is
	port (
		bytesub_0_avalon_streaming_sink_data  : in  std_logic_vector(127 downto 0) := (others => '0'); -- bytesub_0_avalon_streaming_sink.data
		bytesub_0_avalon_streaming_sink_ready : out std_logic;                                         --                                .ready
		bytesub_0_avalon_streaming_sink_valid : in  std_logic                      := '0';             --                                .valid
		clk_clk                               : in  std_logic                      := '0';             --                             clk.clk
		display_0_display_out_data            : out std_logic_vector(7 downto 0);                      --           display_0_display_out.data
		display_1_display_out_data            : out std_logic_vector(7 downto 0);                      --           display_1_display_out.data
		display_2_display_out_data            : out std_logic_vector(7 downto 0);                      --           display_2_display_out.data
		display_3_display_out_data            : out std_logic_vector(7 downto 0);                      --           display_3_display_out.data
		reset_reset_n                         : in  std_logic                      := '0'              --                           reset.reset_n
	);
end entity byteSub_display_sys;

architecture rtl of byteSub_display_sys is
	component byte_sub is
		port (
			clk       : in  std_logic                      := 'X';             -- clk
			reset_n   : in  std_logic                      := 'X';             -- reset_n
			out_valid : out std_logic;                                         -- valid
			out_ready : in  std_logic                      := 'X';             -- ready
			out_data  : out std_logic_vector(127 downto 0);                    -- data
			in_data   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			in_ready  : out std_logic;                                         -- ready
			in_valid  : in  std_logic                      := 'X'              -- valid
		);
	end component byte_sub;

	component display is
		port (
			reset_sink_reset            : in  std_logic                    := 'X';             -- reset
			clock_sink_clk              : in  std_logic                    := 'X';             -- clk
			hex_data                    : out std_logic_vector(7 downto 0);                    -- data
			data_in                     : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			avalon_streaming_sink_ready : out std_logic;                                       -- ready
			avalon_streaming_sink_valid : in  std_logic                    := 'X'              -- valid
		);
	end component display;

	component divider is
		port (
			clk        : in  std_logic                      := 'X';             -- clk
			reset_n    : in  std_logic                      := 'X';             -- reset_n
			in_data    : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			out_data_1 : out std_logic_vector(31 downto 0);                     -- data
			out_data_2 : out std_logic_vector(31 downto 0);                     -- data
			out_data_3 : out std_logic_vector(31 downto 0);                     -- data
			out_data_4 : out std_logic_vector(31 downto 0)                      -- data
		);
	end component divider;

	component byteSub_display_sys_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk   : in  std_logic                      := 'X';             -- clk
			in_rst_0_reset : in  std_logic                      := 'X';             -- reset
			in_0_data      : in  std_logic_vector(127 downto 0) := (others => 'X'); -- data
			in_0_valid     : in  std_logic                      := 'X';             -- valid
			in_0_ready     : out std_logic;                                         -- ready
			out_0_data     : out std_logic_vector(127 downto 0)                     -- data
		);
	end component byteSub_display_sys_avalon_st_adapter;

	component byteSub_display_sys_avalon_st_adapter_001 is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk   : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset : in  std_logic                     := 'X';             -- reset
			in_0_data      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			out_0_data     : out std_logic_vector(7 downto 0);                     -- data
			out_0_valid    : out std_logic;                                        -- valid
			out_0_ready    : in  std_logic                     := 'X'              -- ready
		);
	end component byteSub_display_sys_avalon_st_adapter_001;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal bytesub_0_avalon_streaming_source_valid  : std_logic;                      -- byteSub_0:out_valid -> avalon_st_adapter:in_0_valid
	signal bytesub_0_avalon_streaming_source_data   : std_logic_vector(127 downto 0); -- byteSub_0:out_data -> avalon_st_adapter:in_0_data
	signal bytesub_0_avalon_streaming_source_ready  : std_logic;                      -- avalon_st_adapter:in_0_ready -> byteSub_0:out_ready
	signal avalon_st_adapter_out_0_data             : std_logic_vector(127 downto 0); -- avalon_st_adapter:out_0_data -> divider_0:in_data
	signal divider_0_data_out_1_data                : std_logic_vector(31 downto 0);  -- divider_0:out_data_1 -> avalon_st_adapter_001:in_0_data
	signal avalon_st_adapter_001_out_0_valid        : std_logic;                      -- avalon_st_adapter_001:out_0_valid -> display_0:avalon_streaming_sink_valid
	signal avalon_st_adapter_001_out_0_data         : std_logic_vector(7 downto 0);   -- avalon_st_adapter_001:out_0_data -> display_0:data_in
	signal avalon_st_adapter_001_out_0_ready        : std_logic;                      -- display_0:avalon_streaming_sink_ready -> avalon_st_adapter_001:out_0_ready
	signal divider_0_data_out_2_data                : std_logic_vector(31 downto 0);  -- divider_0:out_data_2 -> avalon_st_adapter_002:in_0_data
	signal avalon_st_adapter_002_out_0_valid        : std_logic;                      -- avalon_st_adapter_002:out_0_valid -> display_1:avalon_streaming_sink_valid
	signal avalon_st_adapter_002_out_0_data         : std_logic_vector(7 downto 0);   -- avalon_st_adapter_002:out_0_data -> display_1:data_in
	signal avalon_st_adapter_002_out_0_ready        : std_logic;                      -- display_1:avalon_streaming_sink_ready -> avalon_st_adapter_002:out_0_ready
	signal divider_0_data_out_3_data                : std_logic_vector(31 downto 0);  -- divider_0:out_data_3 -> avalon_st_adapter_003:in_0_data
	signal avalon_st_adapter_003_out_0_valid        : std_logic;                      -- avalon_st_adapter_003:out_0_valid -> display_2:avalon_streaming_sink_valid
	signal avalon_st_adapter_003_out_0_data         : std_logic_vector(7 downto 0);   -- avalon_st_adapter_003:out_0_data -> display_2:data_in
	signal avalon_st_adapter_003_out_0_ready        : std_logic;                      -- display_2:avalon_streaming_sink_ready -> avalon_st_adapter_003:out_0_ready
	signal divider_0_data_out_4_data                : std_logic_vector(31 downto 0);  -- divider_0:out_data_4 -> avalon_st_adapter_004:in_0_data
	signal avalon_st_adapter_004_out_0_valid        : std_logic;                      -- avalon_st_adapter_004:out_0_valid -> display_3:avalon_streaming_sink_valid
	signal avalon_st_adapter_004_out_0_data         : std_logic_vector(7 downto 0);   -- avalon_st_adapter_004:out_0_data -> display_3:data_in
	signal avalon_st_adapter_004_out_0_ready        : std_logic;                      -- display_3:avalon_streaming_sink_ready -> avalon_st_adapter_004:out_0_ready
	signal rst_controller_reset_out_reset           : std_logic;                      -- rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, avalon_st_adapter_003:in_rst_0_reset, avalon_st_adapter_004:in_rst_0_reset, display_0:reset_sink_reset, display_1:reset_sink_reset, display_2:reset_sink_reset, display_3:reset_sink_reset, rst_controller_reset_out_reset:in]
	signal reset_reset_n_ports_inv                  : std_logic;                      -- reset_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv : std_logic;                      -- rst_controller_reset_out_reset:inv -> [byteSub_0:reset_n, divider_0:reset_n]

begin

	bytesub_0 : component byte_sub
		port map (
			clk       => clk_clk,                                  --                   clock.clk
			reset_n   => rst_controller_reset_out_reset_ports_inv, --                   reset.reset_n
			out_valid => bytesub_0_avalon_streaming_source_valid,  -- avalon_streaming_source.valid
			out_ready => bytesub_0_avalon_streaming_source_ready,  --                        .ready
			out_data  => bytesub_0_avalon_streaming_source_data,   --                        .data
			in_data   => bytesub_0_avalon_streaming_sink_data,     --   avalon_streaming_sink.data
			in_ready  => bytesub_0_avalon_streaming_sink_ready,    --                        .ready
			in_valid  => bytesub_0_avalon_streaming_sink_valid     --                        .valid
		);

	display_0 : component display
		port map (
			reset_sink_reset            => rst_controller_reset_out_reset,    --   reset_sink.reset
			clock_sink_clk              => clk_clk,                           -- clock_sink_1.clk
			hex_data                    => display_0_display_out_data,        --  display_out.data
			data_in                     => avalon_st_adapter_001_out_0_data,  --      data_in.data
			avalon_streaming_sink_ready => avalon_st_adapter_001_out_0_ready, --             .ready
			avalon_streaming_sink_valid => avalon_st_adapter_001_out_0_valid  --             .valid
		);

	display_1 : component display
		port map (
			reset_sink_reset            => rst_controller_reset_out_reset,    --   reset_sink.reset
			clock_sink_clk              => clk_clk,                           -- clock_sink_1.clk
			hex_data                    => display_1_display_out_data,        --  display_out.data
			data_in                     => avalon_st_adapter_002_out_0_data,  --      data_in.data
			avalon_streaming_sink_ready => avalon_st_adapter_002_out_0_ready, --             .ready
			avalon_streaming_sink_valid => avalon_st_adapter_002_out_0_valid  --             .valid
		);

	display_2 : component display
		port map (
			reset_sink_reset            => rst_controller_reset_out_reset,    --   reset_sink.reset
			clock_sink_clk              => clk_clk,                           -- clock_sink_1.clk
			hex_data                    => display_2_display_out_data,        --  display_out.data
			data_in                     => avalon_st_adapter_003_out_0_data,  --      data_in.data
			avalon_streaming_sink_ready => avalon_st_adapter_003_out_0_ready, --             .ready
			avalon_streaming_sink_valid => avalon_st_adapter_003_out_0_valid  --             .valid
		);

	display_3 : component display
		port map (
			reset_sink_reset            => rst_controller_reset_out_reset,    --   reset_sink.reset
			clock_sink_clk              => clk_clk,                           -- clock_sink_1.clk
			hex_data                    => display_3_display_out_data,        --  display_out.data
			data_in                     => avalon_st_adapter_004_out_0_data,  --      data_in.data
			avalon_streaming_sink_ready => avalon_st_adapter_004_out_0_ready, --             .ready
			avalon_streaming_sink_valid => avalon_st_adapter_004_out_0_valid  --             .valid
		);

	divider_0 : component divider
		port map (
			clk        => clk_clk,                                  --      clock.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --      reset.reset_n
			in_data    => avalon_st_adapter_out_0_data,             --    data_in.data
			out_data_1 => divider_0_data_out_1_data,                -- data_out_1.data
			out_data_2 => divider_0_data_out_2_data,                -- data_out_2.data
			out_data_3 => divider_0_data_out_3_data,                -- data_out_3.data
			out_data_4 => divider_0_data_out_4_data                 -- data_out_4.data
		);

	avalon_st_adapter : component byteSub_display_sys_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 0,
			inDataWidth     => 128,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 128,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 0,
			outUseReady     => 0,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => clk_clk,                                 -- in_clk_0.clk
			in_rst_0_reset => rst_controller_reset_out_reset,          -- in_rst_0.reset
			in_0_data      => bytesub_0_avalon_streaming_source_data,  --     in_0.data
			in_0_valid     => bytesub_0_avalon_streaming_source_valid, --         .valid
			in_0_ready     => bytesub_0_avalon_streaming_source_ready, --         .ready
			out_0_data     => avalon_st_adapter_out_0_data             --    out_0.data
		);

	avalon_st_adapter_001 : component byteSub_display_sys_avalon_st_adapter_001
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 0,
			inUseReady      => 0,
			inReadyLatency  => 0,
			outDataWidth    => 8,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => clk_clk,                           -- in_clk_0.clk
			in_rst_0_reset => rst_controller_reset_out_reset,    -- in_rst_0.reset
			in_0_data      => divider_0_data_out_1_data,         --     in_0.data
			out_0_data     => avalon_st_adapter_001_out_0_data,  --    out_0.data
			out_0_valid    => avalon_st_adapter_001_out_0_valid, --         .valid
			out_0_ready    => avalon_st_adapter_001_out_0_ready  --         .ready
		);

	avalon_st_adapter_002 : component byteSub_display_sys_avalon_st_adapter_001
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 0,
			inUseReady      => 0,
			inReadyLatency  => 0,
			outDataWidth    => 8,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => clk_clk,                           -- in_clk_0.clk
			in_rst_0_reset => rst_controller_reset_out_reset,    -- in_rst_0.reset
			in_0_data      => divider_0_data_out_2_data,         --     in_0.data
			out_0_data     => avalon_st_adapter_002_out_0_data,  --    out_0.data
			out_0_valid    => avalon_st_adapter_002_out_0_valid, --         .valid
			out_0_ready    => avalon_st_adapter_002_out_0_ready  --         .ready
		);

	avalon_st_adapter_003 : component byteSub_display_sys_avalon_st_adapter_001
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 0,
			inUseReady      => 0,
			inReadyLatency  => 0,
			outDataWidth    => 8,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => clk_clk,                           -- in_clk_0.clk
			in_rst_0_reset => rst_controller_reset_out_reset,    -- in_rst_0.reset
			in_0_data      => divider_0_data_out_3_data,         --     in_0.data
			out_0_data     => avalon_st_adapter_003_out_0_data,  --    out_0.data
			out_0_valid    => avalon_st_adapter_003_out_0_valid, --         .valid
			out_0_ready    => avalon_st_adapter_003_out_0_ready  --         .ready
		);

	avalon_st_adapter_004 : component byteSub_display_sys_avalon_st_adapter_001
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 0,
			inUseReady      => 0,
			inReadyLatency  => 0,
			outDataWidth    => 8,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => clk_clk,                           -- in_clk_0.clk
			in_rst_0_reset => rst_controller_reset_out_reset,    -- in_rst_0.reset
			in_0_data      => divider_0_data_out_4_data,         --     in_0.data
			out_0_data     => avalon_st_adapter_004_out_0_data,  --    out_0.data
			out_0_valid    => avalon_st_adapter_004_out_0_valid, --         .valid
			out_0_ready    => avalon_st_adapter_004_out_0_ready  --         .ready
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of byteSub_display_sys
