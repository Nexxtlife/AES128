library ieee;
use ieee.std_logic_1164.all;

entity aes_enc is 
	port (
		clk : in std_logic;
		rst : in std_logic;
		key : in std_logic_vector(127 downto 0);
		plaintext : in std_logic_vector(127 downto 0);
		ciphertext : out std_logic_vector(127 downto 0);
		done : out std_logic		
	);
end aes_enc;

architecture behavioral of aes_enc is
	signal inverted_plaintext : std_logic_vector(127 downto 0);
	signal inverted_key : std_logic_vector(127 downto 0);
	signal inverted_cyphertext : std_logic_vector(127 downto 0);
	signal reg_input : std_logic_vector(127 downto 0);
	signal reg_output : std_logic_vector(127 downto 0);
	signal subbox_input : std_logic_vector(127 downto 0);
	signal subbox_output : std_logic_vector(127 downto 0);
	signal shiftrows_output : std_logic_vector(127 downto 0);
	signal mixcol_output : std_logic_vector(127 downto 0);
	signal feedback : std_logic_vector(127 downto 0);
	signal round_key : std_logic_vector(127 downto 0);
	signal round_const : std_logic_vector(7 downto 0);
	signal sel : std_logic;
begin
	inverter_inst_plaintext : entity work.inverter
		port map(
			data_in => plaintext,
			data_out => inverted_plaintext
		);
	inverter_inst_key : entity work.inverter
		port map(
			data_in => key,
			data_out => inverted_key
		);	
	inverter_inst_cyphertext : entity work.inverter
		port map(
			data_in => inverted_cyphertext,
			data_out => ciphertext
		);
	reg_input <= inverted_plaintext when rst = '0' else feedback;
	reg_inst : entity work.reg
		generic map(
			size => 128
		)
		port map(
			clk => clk,
			d   => reg_input,
			q   => reg_output
		);
	-- Encryption body
	add_round_key_inst : entity work.add_round_key
		port map(
			input1 => reg_output,
			input2 => round_key,
			output => subbox_input
		);
	byte_sub_inst : entity work.byte_sub
		port map(
			data_in  => subbox_input,
			data_out => subbox_output
			
		);
	shft_row_inst : entity work.shft_row
		port map(
			data_in  => subbox_output,
			data_out => shiftrows_output
		);
	mix_columns_inst : entity work.mix_column
		port map(
			input_data  => shiftrows_output,
			output_data => mixcol_output
		);
	feedback <= mixcol_output when sel = '0' else shiftrows_output;
	inverted_cyphertext <= subbox_input;	
	-- Controller
	controller_inst : entity work.controller
		port map(
			clk            => clk,
			rst            => rst,
			rconst         => round_const,
			is_final_round => sel,
			done           => done
		);
	-- Keyschedule
	key_schedule_inst : entity work.key_schedule
		port map(
			clk         => clk,
			rst         => rst,
			key         => inverted_key,
			round_const => round_const,
			round_key   => round_key
		);	
end architecture behavioral;