library ieee;
use ieee.std_logic_1164.all;

entity interface_tb is 
end interface_tb;

architecture behavior of interface_tb is
	component interface
		port(
			clk_clk                                   : in  std_logic                      := 'X';             -- clk
			reset_reset_n                             : in  std_logic                      := 'X';             -- reset_n
						
			--interface_0_avalon_master_1_read          : out std_logic;  
			--interface_0_avalon_master_1_waitrequest   : in std_logic;  
			--interface_0_avalon_master_1_address       : out std_logic_vector(16 downto 0);                     -- address
			--interface_0_avalon_master_1_byteenable    : out std_logic_vector(15 downto 0);                     -- byteenable
			--interface_0_avalon_master_1_readdata      : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			
			interface_0_avalon_streaming_source_data  : out std_logic_vector(127 downto 0);                    -- data
			interface_0_avalon_streaming_source_ready : in  std_logic                      := 'X';             -- ready
			interface_0_avalon_streaming_source_valid : out std_logic;                                          -- valid
			
			interface_1_avalon_streaming_sink_data  : in std_logic_vector(127 downto 0);                    -- data
			interface_1_avalon_streaming_sink_ready : out  std_logic;            							  -- ready
			interface_1_avalon_streaming_sink_valid : in std_logic                                          -- valid
	);	
	end component interface;	
	signal clk_tb : std_logic := '0';
	signal rst_tb : std_logic := '0';
	
	signal interface_0_avalon_streaming_source_data_tb : std_logic_vector(127 downto 0);
	signal interface_0_avalon_streaming_source_ready_tb  : std_logic;
	signal interface_0_avalon_streaming_source_valid_tb : std_logic;
			
	signal interface_1_avalon_streaming_sink_data_tb : std_logic_vector(127 downto 0);
	signal interface_1_avalon_streaming_sink_ready_tb  : std_logic;
	signal interface_1_avalon_streaming_sink_valid_tb : std_logic;
	signal plaintext_tb : std_logic_vector(127 downto 0);	
	constant clk_period : time := 10 ns;
	
begin
	interface_inst : interface
		port map(
			clk_clk =>  clk_tb,
			reset_reset_n =>  rst_tb,
								
			interface_0_avalon_streaming_source_data => interface_0_avalon_streaming_source_data_tb,
			interface_0_avalon_streaming_source_ready => interface_0_avalon_streaming_source_ready_tb,
			interface_0_avalon_streaming_source_valid  => interface_0_avalon_streaming_source_valid_tb,
			
			interface_1_avalon_streaming_sink_data => interface_1_avalon_streaming_sink_data_tb,
			interface_1_avalon_streaming_sink_ready => interface_1_avalon_streaming_sink_ready_tb,
			interface_1_avalon_streaming_sink_valid => interface_1_avalon_streaming_sink_valid_tb
	);
	clk_process : process is
	begin
		clk_tb <= '0';
		wait for clk_period/2;
		clk_tb <= '1';
		wait for clk_period/2;
	end process clk_process;
	
	sim_proc : process is
	begin
		report "Testbench started";
		wait until rising_edge(clk_tb) and rst_tb = '0';
		wait until interface_1_avalon_streaming_sink_ready_tb = '1';
		--if(interface_1_avalon_streaming_sink_ready_tb = '1') then
		report "entered if statement";
			interface_1_avalon_streaming_sink_valid_tb <= '1';
			interface_1_avalon_streaming_sink_data_tb <= x"3243f6a8885a308d313198a2e0370734";

			wait for clk_period * 3;
			interface_1_avalon_streaming_sink_valid_tb <='0';
			interface_0_avalon_streaming_source_ready_tb <='1';

			wait for clk_period * 2;
			interface_0_avalon_streaming_source_ready_tb <='1';
		--end if;
	end process sim_proc;
	
	reset_process: process
		variable reset_cycles_count : integer := 2; 
		begin
		rst_tb <= '1';
		while reset_cycles_count >= 0 loop
		  wait until rising_edge(clk_tb);
		  reset_cycles_count := reset_cycles_count - 1;
		end loop;
		rst_tb <= '0';
		--wait for clk_period * 2;
	end process;
	
end architecture behavior;