-- JTAG_AES.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity JTAG_AES is
	port (
		clk_clk         : in std_logic := '0'; --     clk.clk
		reset_n_reset_n : in std_logic := '0'  -- reset_n.reset_n
	);
end entity JTAG_AES;

architecture rtl of JTAG_AES is
	component interface_controller is
		generic (
			INTERFACE_WIDTH      : integer := 32;
			INTERFACE_LENGTH     : natural := 32;
			INTERFACE_ADDR_WIDTH : natural := 5
		);
		port (
			interface_0_avalon_slave_1_read        : in  std_logic                     := 'X';             -- read
			interface_0_avalon_slave_1_write       : in  std_logic                     := 'X';             -- write
			interface_0_avalon_slave_1_waitrequest : out std_logic;                                        -- waitrequest
			interface_0_avalon_slave_1_address     : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			interface_0_avalon_slave_1_byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			interface_0_avalon_slave_1_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			interface_0_avalon_slave_1_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clk_clk                                : in  std_logic                     := 'X';             -- clk
			rst_t                                  : in  std_logic                     := 'X'              -- reset
		);
	end component interface_controller;

	component JTAG_AES_master_0 is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component JTAG_AES_master_0;

	component JTAG_AES_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			AES_0_reset_sink_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			master_0_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			master_0_master_address                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			master_0_master_waitrequest                    : out std_logic;                                        -- waitrequest
			master_0_master_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			master_0_master_read                           : in  std_logic                     := 'X';             -- read
			master_0_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			master_0_master_readdatavalid                  : out std_logic;                                        -- readdatavalid
			master_0_master_write                          : in  std_logic                     := 'X';             -- write
			master_0_master_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			AES_0_interface_0_avalon_slave_1_address       : out std_logic_vector(4 downto 0);                     -- address
			AES_0_interface_0_avalon_slave_1_write         : out std_logic;                                        -- write
			AES_0_interface_0_avalon_slave_1_read          : out std_logic;                                        -- read
			AES_0_interface_0_avalon_slave_1_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			AES_0_interface_0_avalon_slave_1_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			AES_0_interface_0_avalon_slave_1_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			AES_0_interface_0_avalon_slave_1_waitrequest   : in  std_logic                     := 'X'              -- waitrequest
		);
	end component JTAG_AES_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal master_0_master_readdata                                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	signal master_0_master_waitrequest                                    : std_logic;                     -- mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	signal master_0_master_address                                        : std_logic_vector(31 downto 0); -- master_0:master_address -> mm_interconnect_0:master_0_master_address
	signal master_0_master_read                                           : std_logic;                     -- master_0:master_read -> mm_interconnect_0:master_0_master_read
	signal master_0_master_byteenable                                     : std_logic_vector(3 downto 0);  -- master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	signal master_0_master_readdatavalid                                  : std_logic;                     -- mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	signal master_0_master_write                                          : std_logic;                     -- master_0:master_write -> mm_interconnect_0:master_0_master_write
	signal master_0_master_writedata                                      : std_logic_vector(31 downto 0); -- master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	signal mm_interconnect_0_aes_0_interface_0_avalon_slave_1_readdata    : std_logic_vector(31 downto 0); -- AES_0:interface_0_avalon_slave_1_readdata -> mm_interconnect_0:AES_0_interface_0_avalon_slave_1_readdata
	signal mm_interconnect_0_aes_0_interface_0_avalon_slave_1_waitrequest : std_logic;                     -- AES_0:interface_0_avalon_slave_1_waitrequest -> mm_interconnect_0:AES_0_interface_0_avalon_slave_1_waitrequest
	signal mm_interconnect_0_aes_0_interface_0_avalon_slave_1_address     : std_logic_vector(4 downto 0);  -- mm_interconnect_0:AES_0_interface_0_avalon_slave_1_address -> AES_0:interface_0_avalon_slave_1_address
	signal mm_interconnect_0_aes_0_interface_0_avalon_slave_1_read        : std_logic;                     -- mm_interconnect_0:AES_0_interface_0_avalon_slave_1_read -> AES_0:interface_0_avalon_slave_1_read
	signal mm_interconnect_0_aes_0_interface_0_avalon_slave_1_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:AES_0_interface_0_avalon_slave_1_byteenable -> AES_0:interface_0_avalon_slave_1_byteenable
	signal mm_interconnect_0_aes_0_interface_0_avalon_slave_1_write       : std_logic;                     -- mm_interconnect_0:AES_0_interface_0_avalon_slave_1_write -> AES_0:interface_0_avalon_slave_1_write
	signal mm_interconnect_0_aes_0_interface_0_avalon_slave_1_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:AES_0_interface_0_avalon_slave_1_writedata -> AES_0:interface_0_avalon_slave_1_writedata
	signal rst_controller_reset_out_reset                                 : std_logic;                     -- rst_controller:reset_out -> [AES_0:rst_t, mm_interconnect_0:AES_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset]
	signal reset_n_reset_n_ports_inv                                      : std_logic;                     -- reset_n_reset_n:inv -> [master_0:clk_reset_reset, rst_controller:reset_in0]

begin

	aes_0 : component interface_controller
		generic map (
			INTERFACE_WIDTH      => 32,
			INTERFACE_LENGTH     => 32,
			INTERFACE_ADDR_WIDTH => 5
		)
		port map (
			interface_0_avalon_slave_1_read        => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_read,        -- interface_0_avalon_slave_1.read
			interface_0_avalon_slave_1_write       => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_write,       --                           .write
			interface_0_avalon_slave_1_waitrequest => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_waitrequest, --                           .waitrequest
			interface_0_avalon_slave_1_address     => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_address,     --                           .address
			interface_0_avalon_slave_1_byteenable  => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_byteenable,  --                           .byteenable
			interface_0_avalon_slave_1_readdata    => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_readdata,    --                           .readdata
			interface_0_avalon_slave_1_writedata   => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_writedata,   --                           .writedata
			clk_clk                                => clk_clk,                                                        --                 clock_sink.clk
			rst_t                                  => rst_controller_reset_out_reset                                  --                 reset_sink.reset
		);

	master_0 : component JTAG_AES_master_0
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_clk,                       --          clk.clk
			clk_reset_reset      => reset_n_reset_n_ports_inv,     --    clk_reset.reset
			master_address       => master_0_master_address,       --       master.address
			master_readdata      => master_0_master_readdata,      --             .readdata
			master_read          => master_0_master_read,          --             .read
			master_write         => master_0_master_write,         --             .write
			master_writedata     => master_0_master_writedata,     --             .writedata
			master_waitrequest   => master_0_master_waitrequest,   --             .waitrequest
			master_readdatavalid => master_0_master_readdatavalid, --             .readdatavalid
			master_byteenable    => master_0_master_byteenable,    --             .byteenable
			master_reset_reset   => open                           -- master_reset.reset
		);

	mm_interconnect_0 : component JTAG_AES_mm_interconnect_0
		port map (
			clk_0_clk_clk                                  => clk_clk,                                                        --                                clk_0_clk.clk
			AES_0_reset_sink_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                                 --   AES_0_reset_sink_reset_bridge_in_reset.reset
			master_0_clk_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                 -- master_0_clk_reset_reset_bridge_in_reset.reset
			master_0_master_address                        => master_0_master_address,                                        --                          master_0_master.address
			master_0_master_waitrequest                    => master_0_master_waitrequest,                                    --                                         .waitrequest
			master_0_master_byteenable                     => master_0_master_byteenable,                                     --                                         .byteenable
			master_0_master_read                           => master_0_master_read,                                           --                                         .read
			master_0_master_readdata                       => master_0_master_readdata,                                       --                                         .readdata
			master_0_master_readdatavalid                  => master_0_master_readdatavalid,                                  --                                         .readdatavalid
			master_0_master_write                          => master_0_master_write,                                          --                                         .write
			master_0_master_writedata                      => master_0_master_writedata,                                      --                                         .writedata
			AES_0_interface_0_avalon_slave_1_address       => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_address,     --         AES_0_interface_0_avalon_slave_1.address
			AES_0_interface_0_avalon_slave_1_write         => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_write,       --                                         .write
			AES_0_interface_0_avalon_slave_1_read          => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_read,        --                                         .read
			AES_0_interface_0_avalon_slave_1_readdata      => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_readdata,    --                                         .readdata
			AES_0_interface_0_avalon_slave_1_writedata     => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_writedata,   --                                         .writedata
			AES_0_interface_0_avalon_slave_1_byteenable    => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_byteenable,  --                                         .byteenable
			AES_0_interface_0_avalon_slave_1_waitrequest   => mm_interconnect_0_aes_0_interface_0_avalon_slave_1_waitrequest  --                                         .waitrequest
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_n_reset_n_ports_inv,      -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_n_reset_n_ports_inv <= not reset_n_reset_n;

end architecture rtl; -- of JTAG_AES
